library verilog;
use verilog.vl_types.all;
entity TesteMemoriaInst_vlg_vec_tst is
end TesteMemoriaInst_vlg_vec_tst;
