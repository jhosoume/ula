library verilog;
use verilog.vl_types.all;
entity TesteCounter_vlg_vec_tst is
end TesteCounter_vlg_vec_tst;
