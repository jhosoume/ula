library verilog;
use verilog.vl_types.all;
entity ZeroExtensor_vlg_vec_tst is
end ZeroExtensor_vlg_vec_tst;
