library verilog;
use verilog.vl_types.all;
entity TesteAdder32_vlg_vec_tst is
end TesteAdder32_vlg_vec_tst;
