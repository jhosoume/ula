library verilog;
use verilog.vl_types.all;
entity MemoriaInstrucoesFinal_vlg_vec_tst is
end MemoriaInstrucoesFinal_vlg_vec_tst;
