library verilog;
use verilog.vl_types.all;
entity MemoryControl_vlg_vec_tst is
end MemoryControl_vlg_vec_tst;
