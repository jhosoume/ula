    Mac OS X            	   2   �      �                                      ATTR       �   �   S                  �   S  com.dropbox.attributes   x��VJ)�/Hʯ�O��I�L���ON�Q�R�V�ML����%����RK�%�B��D7S�� ����2�$˰|/G[[���Z �,J