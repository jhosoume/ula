library verilog;
use verilog.vl_types.all;
entity SinalExtensor_vlg_vec_tst is
end SinalExtensor_vlg_vec_tst;
