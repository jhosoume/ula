library verilog;
use verilog.vl_types.all;
entity TesteMUX2_vlg_check_tst is
    port(
        Y               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end TesteMUX2_vlg_check_tst;
