library verilog;
use verilog.vl_types.all;
entity NovoBancoDeRegistradores_vlg_vec_tst is
end NovoBancoDeRegistradores_vlg_vec_tst;
