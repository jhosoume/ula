library verilog;
use verilog.vl_types.all;
entity FreqDiv_vlg_check_tst is
    port(
        Div2            : in     vl_logic;
        Div4            : in     vl_logic;
        Div8            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end FreqDiv_vlg_check_tst;
