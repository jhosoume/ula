library verilog;
use verilog.vl_types.all;
entity TesteShiftRegister_vlg_vec_tst is
end TesteShiftRegister_vlg_vec_tst;
