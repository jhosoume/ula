library verilog;
use verilog.vl_types.all;
entity TesteMainULA_vlg_vec_tst is
end TesteMainULA_vlg_vec_tst;
