library verilog;
use verilog.vl_types.all;
entity FreqDiv_vlg_vec_tst is
end FreqDiv_vlg_vec_tst;
