library verilog;
use verilog.vl_types.all;
entity SumSub_vlg_vec_tst is
end SumSub_vlg_vec_tst;
