library verilog;
use verilog.vl_types.all;
entity Mult_vlg_vec_tst is
end Mult_vlg_vec_tst;
