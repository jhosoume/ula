library verilog;
use verilog.vl_types.all;
entity TesteFioBUS_vlg_vec_tst is
end TesteFioBUS_vlg_vec_tst;
