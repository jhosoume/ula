library verilog;
use verilog.vl_types.all;
entity LoadUpperImmediate_vlg_vec_tst is
end LoadUpperImmediate_vlg_vec_tst;
