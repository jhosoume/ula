library verilog;
use verilog.vl_types.all;
entity GetAddrs_vlg_vec_tst is
end GetAddrs_vlg_vec_tst;
