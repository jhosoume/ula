library verilog;
use verilog.vl_types.all;
entity TesteMUX2_vlg_vec_tst is
end TesteMUX2_vlg_vec_tst;
