library verilog;
use verilog.vl_types.all;
entity TesteShift2BitsLeft_vlg_vec_tst is
end TesteShift2BitsLeft_vlg_vec_tst;
