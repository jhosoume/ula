library verilog;
use verilog.vl_types.all;
entity teste_ula_1bit_vlg_vec_tst is
end teste_ula_1bit_vlg_vec_tst;
