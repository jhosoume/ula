library verilog;
use verilog.vl_types.all;
entity TesteRegister_vlg_vec_tst is
end TesteRegister_vlg_vec_tst;
