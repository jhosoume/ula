library verilog;
use verilog.vl_types.all;
entity Keyboard_vlg_vec_tst is
end Keyboard_vlg_vec_tst;
