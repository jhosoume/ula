library verilog;
use verilog.vl_types.all;
entity NewMemoryControl_vlg_vec_tst is
end NewMemoryControl_vlg_vec_tst;
