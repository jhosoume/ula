library verilog;
use verilog.vl_types.all;
entity ZeroExtensor_Shamt_vlg_vec_tst is
end ZeroExtensor_Shamt_vlg_vec_tst;
