    Mac OS X            	   2   �      �                                      ATTR       �   �   S                  �   S  com.dropbox.attributes   x��VJ)�/Hʯ�O��I�L���ON�Q�R�V�ML����%����RK���_��
_߀tm�|o�䤈�t[[���Z Ϋ�