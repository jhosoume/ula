library verilog;
use verilog.vl_types.all;
entity TesteAdd4_vlg_vec_tst is
end TesteAdd4_vlg_vec_tst;
