library verilog;
use verilog.vl_types.all;
entity TesteAdd4_vlg_check_tst is
    port(
        R               : in     vl_logic_vector(31 downto 0);
        sampler_rx      : in     vl_logic
    );
end TesteAdd4_vlg_check_tst;
