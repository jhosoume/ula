library verilog;
use verilog.vl_types.all;
entity ShiftRegister32_vlg_vec_tst is
end ShiftRegister32_vlg_vec_tst;
