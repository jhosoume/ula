library verilog;
use verilog.vl_types.all;
entity Keyboard_vlg_check_tst is
    port(
        KEYINPUT        : in     vl_logic_vector(3 downto 0);
        OUTPUT          : in     vl_logic_vector(7 downto 0);
        sampler_rx      : in     vl_logic
    );
end Keyboard_vlg_check_tst;
