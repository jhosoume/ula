library verilog;
use verilog.vl_types.all;
entity TesteMemoryControl_vlg_vec_tst is
end TesteMemoryControl_vlg_vec_tst;
