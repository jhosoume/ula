library verilog;
use verilog.vl_types.all;
entity TesteInstructionMemory_vlg_vec_tst is
end TesteInstructionMemory_vlg_vec_tst;
