library verilog;
use verilog.vl_types.all;
entity RingCounter_vlg_vec_tst is
end RingCounter_vlg_vec_tst;
