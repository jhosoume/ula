library verilog;
use verilog.vl_types.all;
entity testeMUXBUS_vlg_vec_tst is
end testeMUXBUS_vlg_vec_tst;
