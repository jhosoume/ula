library verilog;
use verilog.vl_types.all;
entity teste_fios_vlg_vec_tst is
end teste_fios_vlg_vec_tst;
