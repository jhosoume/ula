library verilog;
use verilog.vl_types.all;
entity MemoriaDados_vlg_vec_tst is
end MemoriaDados_vlg_vec_tst;
