library verilog;
use verilog.vl_types.all;
entity SignalExtensor_vlg_vec_tst is
end SignalExtensor_vlg_vec_tst;
