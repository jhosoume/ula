library verilog;
use verilog.vl_types.all;
entity Shift2BitsLeft_vlg_vec_tst is
end Shift2BitsLeft_vlg_vec_tst;
